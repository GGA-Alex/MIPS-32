module shoftLeft2(
	input [25:0] entrada,
	output [27:0] salida
);

assign salida = entrada << 2;

endmodule

